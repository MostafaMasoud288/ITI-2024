module instruction_memory
(
input [7:0] A,
output [31:0] RD
);
reg [31:0] ROM [0:255];
integer i;
initial
begin

ROM[0]=32'h00500113;
ROM[1]=32'h00C00193;
ROM[2]=32'hFF718393;
ROM[3]=32'h0023E233;
ROM[4]=32'h0041F2B3;
ROM[5]=32'h004282B3;
ROM[6]=32'h02728863;
ROM[7]=32'h0041A233;
ROM[8]=32'h00020463;
ROM[9]=32'h00000293;
ROM[10]=32'h0023A233;
ROM[11]=32'h005203B3;
ROM[12]=32'h402383B3;
ROM[13]=32'h0471AA23;
ROM[14]=32'h06002103;
ROM[15]=32'h005104B3;
ROM[16]=32'h008001EF;
ROM[17]=32'h00100113;
ROM[18]=32'h00910133;
ROM[19]=32'h0221A023;
ROM[20]=32'h00210063;
for(i=21;i<256;i=i+1)
ROM[i]=32'h0;/*
ROM[0]  = 32'b00000000101000000000000010010011;  // addi x1, x0, 10
ROM[1]  = 32'b00000001010000000000000100010011;  // addi x2, x0, 20
ROM[2]  = 32'b00000010100000000000000110010011;  // addi x3, x0, 40
ROM[3]  = 32'b00000101000000000000001000010011;  // addi x4, x0, 80
ROM[4]  = 32'b00001010000000000000001010010011;  // addi x5, x0, 160
ROM[5]  = 32'b00000000000100000010000000100011;  // sw x1, 0(x0)
ROM[6]  = 32'b00000000001000000010001000100011;  // sw x2, 4(x0)
ROM[7]  = 32'b00000000001100000010010000100011;  // sw x3, 8(x0)
ROM[8]  = 32'b00000000010000000010011000100011;  // sw x4, 12(x0)
ROM[9]  = 32'b00000000010100000010011000100011;  // sw x5, 12(x0)
ROM[10]  = 32'b00000000000000000010010100000011;  // lw x10, 0(x0)
ROM[11] = 32'b00000000010000000010010110000011;  // lw x11, 4(x0)
ROM[12] = 32'b00000000100000000010011000000011;  // lw x12, 8(x0)
ROM[13] = 32'b00000000110000000010011010000011;  // lw x13, 12(x0)
ROM[14] = 32'b00000000010000000010011000100011;  //�sw�x4,�12(x0)
for(i=15;i<256;i=i+1)
ROM[i]=32'h0;*/
end
assign RD = ROM[A];
endmodule